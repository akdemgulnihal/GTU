magic
tech scmos
timestamp 1706367479
<< nwell >>
rect -25 -6 -1 16
<< ntransistor >>
rect -14 -20 -12 -16
<< ptransistor >>
rect -14 0 -12 4
<< ndiffusion >>
rect -15 -20 -14 -16
rect -12 -20 -11 -16
<< pdiffusion >>
rect -15 0 -14 4
rect -12 0 -11 4
<< ndcontact >>
rect -19 -20 -15 -16
rect -11 -20 -7 -16
<< pdcontact >>
rect -19 0 -15 4
rect -11 0 -7 4
<< psubstratepcontact >>
rect -17 -29 -7 -25
<< nsubstratencontact >>
rect -18 9 -8 13
<< polysilicon >>
rect -14 4 -12 7
rect -14 -6 -12 0
rect -16 -10 -12 -6
rect -14 -16 -12 -10
rect -14 -23 -12 -20
<< polycontact >>
rect -20 -10 -16 -6
<< metal1 >>
rect -23 13 -3 14
rect -23 9 -18 13
rect -8 9 -3 13
rect -23 8 -3 9
rect -19 4 -15 8
rect -11 -6 -7 0
rect -24 -10 -20 -6
rect -11 -10 -3 -6
rect -11 -16 -7 -10
rect -19 -24 -15 -20
rect -23 -25 -3 -24
rect -23 -29 -17 -25
rect -7 -29 -3 -25
rect -23 -30 -3 -29
<< labels >>
rlabel metal1 -21 -26 -21 -26 2 Gnd
rlabel metal1 -22 12 -22 12 4 Vdd
<< end >>
