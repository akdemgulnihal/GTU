magic
tech scmos
timestamp 1703861445
<< nwell >>
rect -17 -3 33 19
<< ntransistor >>
rect -6 -28 -4 -24
rect 1 -28 3 -24
rect 10 -28 12 -24
rect 18 -28 20 -24
<< ptransistor >>
rect -6 3 -4 7
rect 1 3 3 7
rect 10 3 12 7
rect 18 3 20 7
<< ndiffusion >>
rect -7 -28 -6 -24
rect -4 -28 1 -24
rect 3 -28 4 -24
rect 8 -28 10 -24
rect 12 -28 18 -24
rect 20 -28 21 -24
<< pdiffusion >>
rect -7 3 -6 7
rect -4 3 1 7
rect 3 3 4 7
rect 8 3 10 7
rect 12 3 13 7
rect 17 3 18 7
rect 20 3 21 7
<< ndcontact >>
rect -11 -28 -7 -24
rect 4 -28 8 -24
rect 21 -28 25 -24
<< pdcontact >>
rect -11 3 -7 7
rect 4 3 8 7
rect 13 3 17 7
rect 21 3 25 7
<< psubstratepcontact >>
rect -11 -37 -7 -33
rect 19 -37 23 -33
<< nsubstratencontact >>
rect -12 12 -8 16
rect -4 12 0 16
<< polysilicon >>
rect -6 8 -4 10
rect 1 8 3 10
rect 10 8 12 10
rect 18 8 20 10
rect -6 -8 -4 3
rect 1 -7 3 3
rect 10 -8 12 3
rect 18 -8 20 3
rect -6 -24 -4 -13
rect 1 -24 3 -12
rect 10 -24 12 -13
rect 18 -24 20 -13
rect -6 -31 -4 -28
rect 1 -31 3 -28
rect 10 -31 12 -28
rect 18 -31 20 -28
<< polycontact >>
rect -9 -13 -4 -8
rect 0 -12 5 -7
rect 9 -13 14 -8
rect 18 -13 23 -8
<< polypplus >>
rect -6 7 -4 8
rect 1 7 3 8
rect 10 7 12 8
rect 18 7 20 8
<< metal1 >>
rect -12 16 0 17
rect -8 12 -4 16
rect -12 11 0 12
rect -3 4 0 11
rect 4 11 25 14
rect 4 7 8 11
rect 21 7 25 11
rect -11 1 -7 3
rect 4 1 8 3
rect -11 -2 8 1
rect 13 0 17 3
rect 13 -3 30 0
rect 27 -18 30 -3
rect -11 -21 30 -18
rect -11 -24 -7 -21
rect 21 -24 25 -21
rect 4 -32 8 -28
rect -12 -33 24 -32
rect -12 -37 -11 -33
rect -7 -37 19 -33
rect 23 -37 24 -33
rect -12 -38 24 -37
<< labels >>
rlabel metal1 5 -34 5 -34 1 Gnd
rlabel metal1 -6 14 -6 14 5 VDD
<< end >>
