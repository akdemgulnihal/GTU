magic
tech scmos
timestamp 1702478130
<< nwell >>
rect -219 0 -83 32
rect -7 4 129 36
rect 300 2 436 34
rect 512 6 648 38
<< ntransistor >>
rect 5 -19 7 -15
rect 21 -19 23 -15
rect 29 -19 31 -15
rect 37 -19 39 -15
rect 45 -19 47 -15
rect 51 -19 53 -15
rect 59 -19 61 -15
rect 67 -19 69 -15
rect 75 -19 77 -15
rect 83 -19 85 -15
rect 93 -19 95 -15
rect 99 -19 101 -15
rect 105 -19 107 -15
rect 113 -19 115 -15
rect 524 -17 526 -13
rect 540 -17 542 -13
rect 548 -17 550 -13
rect 556 -17 558 -13
rect 564 -17 566 -13
rect 570 -17 572 -13
rect 578 -17 580 -13
rect 586 -17 588 -13
rect 594 -17 596 -13
rect 602 -17 604 -13
rect 612 -17 614 -13
rect 618 -17 620 -13
rect 624 -17 626 -13
rect 632 -17 634 -13
rect -207 -23 -205 -19
rect -191 -23 -189 -19
rect -183 -23 -181 -19
rect -175 -23 -173 -19
rect -167 -23 -165 -19
rect -161 -23 -159 -19
rect -153 -23 -151 -19
rect -145 -23 -143 -19
rect -137 -23 -135 -19
rect -129 -23 -127 -19
rect -119 -23 -117 -19
rect -113 -23 -111 -19
rect -107 -23 -105 -19
rect -99 -23 -97 -19
rect 312 -21 314 -17
rect 328 -21 330 -17
rect 336 -21 338 -17
rect 344 -21 346 -17
rect 352 -21 354 -17
rect 358 -21 360 -17
rect 366 -21 368 -17
rect 374 -21 376 -17
rect 382 -21 384 -17
rect 390 -21 392 -17
rect 400 -21 402 -17
rect 406 -21 408 -17
rect 412 -21 414 -17
rect 420 -21 422 -17
<< ptransistor >>
rect 5 12 7 16
rect 21 12 23 16
rect 29 12 31 16
rect 37 12 39 16
rect 45 12 47 16
rect 51 12 53 16
rect 59 12 61 16
rect 67 12 69 16
rect 75 12 77 16
rect 83 12 85 16
rect 93 12 95 16
rect 99 12 101 16
rect 105 12 107 16
rect 113 12 115 16
rect 524 14 526 18
rect 540 14 542 18
rect 548 14 550 18
rect 556 14 558 18
rect 564 14 566 18
rect 570 14 572 18
rect 578 14 580 18
rect 586 14 588 18
rect 594 14 596 18
rect 602 14 604 18
rect 612 14 614 18
rect 618 14 620 18
rect 624 14 626 18
rect 632 14 634 18
rect -207 8 -205 12
rect -191 8 -189 12
rect -183 8 -181 12
rect -175 8 -173 12
rect -167 8 -165 12
rect -161 8 -159 12
rect -153 8 -151 12
rect -145 8 -143 12
rect -137 8 -135 12
rect -129 8 -127 12
rect -119 8 -117 12
rect -113 8 -111 12
rect -107 8 -105 12
rect -99 8 -97 12
rect 312 10 314 14
rect 328 10 330 14
rect 336 10 338 14
rect 344 10 346 14
rect 352 10 354 14
rect 358 10 360 14
rect 366 10 368 14
rect 374 10 376 14
rect 382 10 384 14
rect 390 10 392 14
rect 400 10 402 14
rect 406 10 408 14
rect 412 10 414 14
rect 420 10 422 14
<< ndiffusion >>
rect 4 -19 5 -15
rect 7 -19 8 -15
rect 20 -19 21 -15
rect 23 -19 24 -15
rect 28 -19 29 -15
rect 31 -19 32 -15
rect 36 -19 37 -15
rect 39 -19 40 -15
rect 44 -19 45 -15
rect 47 -19 51 -15
rect 53 -19 54 -15
rect 58 -19 59 -15
rect 61 -19 62 -15
rect 66 -19 67 -15
rect 69 -19 70 -15
rect 74 -19 75 -15
rect 77 -19 78 -15
rect 82 -19 83 -15
rect 85 -19 88 -15
rect 92 -19 93 -15
rect 95 -19 99 -15
rect 101 -19 105 -15
rect 107 -19 108 -15
rect 112 -19 113 -15
rect 115 -19 119 -15
rect 523 -17 524 -13
rect 526 -17 527 -13
rect 539 -17 540 -13
rect 542 -17 543 -13
rect 547 -17 548 -13
rect 550 -17 551 -13
rect 555 -17 556 -13
rect 558 -17 559 -13
rect 563 -17 564 -13
rect 566 -17 570 -13
rect 572 -17 573 -13
rect 577 -17 578 -13
rect 580 -17 581 -13
rect 585 -17 586 -13
rect 588 -17 589 -13
rect 593 -17 594 -13
rect 596 -17 597 -13
rect 601 -17 602 -13
rect 604 -17 607 -13
rect 611 -17 612 -13
rect 614 -17 618 -13
rect 620 -17 624 -13
rect 626 -17 627 -13
rect 631 -17 632 -13
rect 634 -17 638 -13
rect -208 -23 -207 -19
rect -205 -23 -204 -19
rect -192 -23 -191 -19
rect -189 -23 -188 -19
rect -184 -23 -183 -19
rect -181 -23 -180 -19
rect -176 -23 -175 -19
rect -173 -23 -172 -19
rect -168 -23 -167 -19
rect -165 -23 -161 -19
rect -159 -23 -158 -19
rect -154 -23 -153 -19
rect -151 -23 -150 -19
rect -146 -23 -145 -19
rect -143 -23 -142 -19
rect -138 -23 -137 -19
rect -135 -23 -134 -19
rect -130 -23 -129 -19
rect -127 -23 -124 -19
rect -120 -23 -119 -19
rect -117 -23 -113 -19
rect -111 -23 -107 -19
rect -105 -23 -104 -19
rect -100 -23 -99 -19
rect -97 -23 -93 -19
rect 311 -21 312 -17
rect 314 -21 315 -17
rect 327 -21 328 -17
rect 330 -21 331 -17
rect 335 -21 336 -17
rect 338 -21 339 -17
rect 343 -21 344 -17
rect 346 -21 347 -17
rect 351 -21 352 -17
rect 354 -21 358 -17
rect 360 -21 361 -17
rect 365 -21 366 -17
rect 368 -21 369 -17
rect 373 -21 374 -17
rect 376 -21 377 -17
rect 381 -21 382 -17
rect 384 -21 385 -17
rect 389 -21 390 -17
rect 392 -21 395 -17
rect 399 -21 400 -17
rect 402 -21 406 -17
rect 408 -21 412 -17
rect 414 -21 415 -17
rect 419 -21 420 -17
rect 422 -21 426 -17
<< pdiffusion >>
rect 4 12 5 16
rect 7 12 8 16
rect 20 12 21 16
rect 23 12 24 16
rect 28 12 29 16
rect 31 12 32 16
rect 36 12 37 16
rect 39 12 40 16
rect 44 12 45 16
rect 47 12 51 16
rect 53 12 54 16
rect 58 12 59 16
rect 61 12 62 16
rect 66 12 67 16
rect 69 12 70 16
rect 74 12 75 16
rect 77 12 78 16
rect 82 12 83 16
rect 85 12 88 16
rect 92 12 93 16
rect 95 12 99 16
rect 101 12 105 16
rect 107 12 108 16
rect 112 12 113 16
rect 115 12 119 16
rect 523 14 524 18
rect 526 14 527 18
rect 539 14 540 18
rect 542 14 543 18
rect 547 14 548 18
rect 550 14 551 18
rect 555 14 556 18
rect 558 14 559 18
rect 563 14 564 18
rect 566 14 570 18
rect 572 14 573 18
rect 577 14 578 18
rect 580 14 581 18
rect 585 14 586 18
rect 588 14 589 18
rect 593 14 594 18
rect 596 14 597 18
rect 601 14 602 18
rect 604 14 607 18
rect 611 14 612 18
rect 614 14 618 18
rect 620 14 624 18
rect 626 14 627 18
rect 631 14 632 18
rect 634 14 638 18
rect -208 8 -207 12
rect -205 8 -204 12
rect -192 8 -191 12
rect -189 8 -188 12
rect -184 8 -183 12
rect -181 8 -180 12
rect -176 8 -175 12
rect -173 8 -172 12
rect -168 8 -167 12
rect -165 8 -161 12
rect -159 8 -158 12
rect -154 8 -153 12
rect -151 8 -150 12
rect -146 8 -145 12
rect -143 8 -142 12
rect -138 8 -137 12
rect -135 8 -134 12
rect -130 8 -129 12
rect -127 8 -124 12
rect -120 8 -119 12
rect -117 8 -113 12
rect -111 8 -107 12
rect -105 8 -104 12
rect -100 8 -99 12
rect -97 8 -93 12
rect 311 10 312 14
rect 314 10 315 14
rect 327 10 328 14
rect 330 10 331 14
rect 335 10 336 14
rect 338 10 339 14
rect 343 10 344 14
rect 346 10 347 14
rect 351 10 352 14
rect 354 10 358 14
rect 360 10 361 14
rect 365 10 366 14
rect 368 10 369 14
rect 373 10 374 14
rect 376 10 377 14
rect 381 10 382 14
rect 384 10 385 14
rect 389 10 390 14
rect 392 10 395 14
rect 399 10 400 14
rect 402 10 406 14
rect 408 10 412 14
rect 414 10 415 14
rect 419 10 420 14
rect 422 10 426 14
<< ndcontact >>
rect 0 -19 4 -15
rect 8 -19 12 -15
rect 16 -19 20 -15
rect 24 -19 28 -15
rect 32 -19 36 -15
rect 40 -19 44 -15
rect 54 -19 58 -15
rect 62 -19 66 -15
rect 70 -19 74 -15
rect 78 -19 82 -15
rect 88 -19 92 -15
rect 108 -19 112 -15
rect 119 -19 123 -15
rect 519 -17 523 -13
rect 527 -17 531 -13
rect 535 -17 539 -13
rect 543 -17 547 -13
rect 551 -17 555 -13
rect 559 -17 563 -13
rect 573 -17 577 -13
rect 581 -17 585 -13
rect 589 -17 593 -13
rect 597 -17 601 -13
rect 607 -17 611 -13
rect 627 -17 631 -13
rect 638 -17 642 -13
rect -212 -23 -208 -19
rect -204 -23 -200 -19
rect -196 -23 -192 -19
rect -188 -23 -184 -19
rect -180 -23 -176 -19
rect -172 -23 -168 -19
rect -158 -23 -154 -19
rect -150 -23 -146 -19
rect -142 -23 -138 -19
rect -134 -23 -130 -19
rect -124 -23 -120 -19
rect -104 -23 -100 -19
rect -93 -23 -89 -19
rect 307 -21 311 -17
rect 315 -21 319 -17
rect 323 -21 327 -17
rect 331 -21 335 -17
rect 339 -21 343 -17
rect 347 -21 351 -17
rect 361 -21 365 -17
rect 369 -21 373 -17
rect 377 -21 381 -17
rect 385 -21 389 -17
rect 395 -21 399 -17
rect 415 -21 419 -17
rect 426 -21 430 -17
<< pdcontact >>
rect 0 12 4 16
rect 8 12 12 16
rect 16 12 20 16
rect 24 12 28 16
rect 32 12 36 16
rect 40 12 44 16
rect 54 12 58 16
rect 62 12 66 16
rect 70 12 74 16
rect 78 12 82 16
rect 88 12 92 16
rect 108 12 112 16
rect 119 12 123 16
rect 519 14 523 18
rect 527 14 531 18
rect 535 14 539 18
rect 543 14 547 18
rect 551 14 555 18
rect 559 14 563 18
rect 573 14 577 18
rect 581 14 585 18
rect 589 14 593 18
rect 597 14 601 18
rect 607 14 611 18
rect 627 14 631 18
rect 638 14 642 18
rect -212 8 -208 12
rect -204 8 -200 12
rect -196 8 -192 12
rect -188 8 -184 12
rect -180 8 -176 12
rect -172 8 -168 12
rect -158 8 -154 12
rect -150 8 -146 12
rect -142 8 -138 12
rect -134 8 -130 12
rect -124 8 -120 12
rect -104 8 -100 12
rect -93 8 -89 12
rect 307 10 311 14
rect 315 10 319 14
rect 323 10 327 14
rect 331 10 335 14
rect 339 10 343 14
rect 347 10 351 14
rect 361 10 365 14
rect 369 10 373 14
rect 377 10 381 14
rect 385 10 389 14
rect 395 10 399 14
rect 415 10 419 14
rect 426 10 430 14
<< psubstratepcontact >>
rect -3 -38 1 -34
rect 5 -38 9 -34
rect 516 -36 520 -32
rect 524 -36 528 -32
rect -215 -42 -211 -38
rect -207 -42 -203 -38
rect 304 -40 308 -36
rect 312 -40 316 -36
<< nsubstratencontact >>
rect -215 19 -211 23
rect -207 19 -203 23
rect -3 23 1 27
rect 5 23 9 27
rect 304 21 308 25
rect 312 21 316 25
rect 516 25 520 29
rect 524 25 528 29
<< polysilicon >>
rect 41 35 107 37
rect 560 37 626 39
rect -171 31 -105 33
rect -207 12 -205 15
rect -191 12 -189 23
rect -183 12 -181 23
rect -175 12 -173 30
rect -167 12 -165 15
rect -161 12 -159 23
rect -153 12 -151 15
rect -145 12 -143 23
rect -137 12 -135 31
rect -129 12 -127 15
rect -119 12 -117 23
rect -113 12 -111 15
rect -107 12 -105 31
rect 5 16 7 19
rect 21 16 23 27
rect 29 16 31 27
rect 37 16 39 34
rect 45 16 47 19
rect 51 16 53 27
rect 59 16 61 19
rect 67 16 69 27
rect 75 16 77 35
rect 83 16 85 19
rect 93 16 95 27
rect 99 16 101 19
rect 105 16 107 35
rect 348 33 414 35
rect 113 16 115 19
rect -99 12 -97 15
rect 312 14 314 17
rect 328 14 330 25
rect 336 14 338 25
rect 344 14 346 32
rect 352 14 354 17
rect 358 14 360 25
rect 366 14 368 17
rect 374 14 376 25
rect 382 14 384 33
rect 390 14 392 17
rect 400 14 402 25
rect 406 14 408 17
rect 412 14 414 33
rect 524 18 526 21
rect 540 18 542 29
rect 548 18 550 29
rect 556 18 558 36
rect 564 18 566 21
rect 570 18 572 29
rect 578 18 580 21
rect 586 18 588 29
rect 594 18 596 37
rect 602 18 604 21
rect 612 18 614 29
rect 618 18 620 21
rect 624 18 626 37
rect 632 18 634 21
rect 420 14 422 17
rect -207 -19 -205 8
rect -191 -19 -189 8
rect -183 -19 -181 8
rect -175 -19 -173 8
rect -167 -19 -165 8
rect -161 -19 -159 8
rect -153 -19 -151 8
rect -145 -19 -143 8
rect -137 -19 -135 8
rect -129 -3 -127 8
rect -129 -19 -127 -7
rect -119 -19 -117 8
rect -113 -19 -111 8
rect -107 -19 -105 8
rect -99 -3 -97 8
rect -99 -19 -97 -7
rect 5 -15 7 12
rect 21 -15 23 12
rect 29 -15 31 12
rect 37 -15 39 12
rect 45 -15 47 12
rect 51 -15 53 12
rect 59 -15 61 12
rect 67 -15 69 12
rect 75 -15 77 12
rect 83 1 85 12
rect 83 -15 85 -3
rect 93 -15 95 12
rect 99 -15 101 12
rect 105 -15 107 12
rect 113 1 115 12
rect 113 -15 115 -3
rect 312 -17 314 10
rect 328 -17 330 10
rect 336 -17 338 10
rect 344 -17 346 10
rect 352 -17 354 10
rect 358 -17 360 10
rect 366 -17 368 10
rect 374 -17 376 10
rect 382 -17 384 10
rect 390 -1 392 10
rect 390 -17 392 -5
rect 400 -17 402 10
rect 406 -17 408 10
rect 412 -17 414 10
rect 420 -1 422 10
rect 420 -17 422 -5
rect 524 -13 526 14
rect 540 -13 542 14
rect 548 -13 550 14
rect 556 -13 558 14
rect 564 -13 566 14
rect 570 -13 572 14
rect 578 -13 580 14
rect 586 -13 588 14
rect 594 -13 596 14
rect 602 3 604 14
rect 602 -13 604 -1
rect 612 -13 614 14
rect 618 -13 620 14
rect 624 -13 626 14
rect 632 3 634 14
rect 632 -13 634 -1
rect 5 -22 7 -19
rect -207 -26 -205 -23
rect -191 -32 -189 -23
rect -183 -26 -181 -23
rect -175 -26 -173 -23
rect -167 -32 -165 -23
rect -161 -26 -159 -23
rect -153 -32 -151 -23
rect -145 -26 -143 -23
rect -137 -26 -135 -23
rect -129 -26 -127 -23
rect -119 -26 -117 -23
rect -113 -32 -111 -23
rect -107 -26 -105 -23
rect -99 -26 -97 -23
rect 21 -28 23 -19
rect 29 -22 31 -19
rect 37 -22 39 -19
rect 45 -28 47 -19
rect 51 -22 53 -19
rect 59 -28 61 -19
rect 67 -22 69 -19
rect 75 -22 77 -19
rect 83 -22 85 -19
rect 93 -22 95 -19
rect 99 -28 101 -19
rect 105 -22 107 -19
rect 113 -22 115 -19
rect 524 -20 526 -17
rect 312 -24 314 -21
rect 21 -30 101 -28
rect 328 -30 330 -21
rect 336 -24 338 -21
rect 344 -24 346 -21
rect 352 -30 354 -21
rect 358 -24 360 -21
rect 366 -30 368 -21
rect 374 -24 376 -21
rect 382 -24 384 -21
rect 390 -24 392 -21
rect 400 -24 402 -21
rect 406 -30 408 -21
rect 412 -24 414 -21
rect 420 -24 422 -21
rect 540 -26 542 -17
rect 548 -20 550 -17
rect 556 -20 558 -17
rect 564 -26 566 -17
rect 570 -20 572 -17
rect 578 -26 580 -17
rect 586 -20 588 -17
rect 594 -20 596 -17
rect 602 -20 604 -17
rect 612 -20 614 -17
rect 618 -26 620 -17
rect 624 -20 626 -17
rect 632 -20 634 -17
rect 540 -28 620 -26
rect 328 -32 408 -30
rect -191 -34 -111 -32
<< polycontact >>
rect 37 34 41 38
rect 556 36 560 40
rect -175 30 -171 34
rect -192 23 -188 27
rect -183 23 -179 27
rect -162 23 -158 27
rect -146 23 -142 27
rect -120 23 -116 27
rect 20 27 24 31
rect 29 27 33 31
rect 50 27 54 31
rect 66 27 70 31
rect 92 27 96 31
rect 344 32 348 36
rect 327 25 331 29
rect 336 25 340 29
rect 357 25 361 29
rect 373 25 377 29
rect 399 25 403 29
rect 539 29 543 33
rect 548 29 552 33
rect 569 29 573 33
rect 585 29 589 33
rect 611 29 615 33
rect -205 -7 -201 -3
rect -131 -7 -127 -3
rect -100 -7 -96 -3
rect 7 -3 11 1
rect 81 -3 85 1
rect 112 -3 116 1
rect 314 -5 318 -1
rect 388 -5 392 -1
rect 419 -5 423 -1
rect 526 -1 530 3
rect 600 -1 604 3
rect 631 -1 635 3
<< metal1 >>
rect 344 47 462 51
rect -175 37 -56 42
rect -175 34 -171 37
rect -216 23 -202 24
rect -179 23 -162 27
rect -158 23 -146 27
rect -142 23 -120 27
rect -216 19 -215 23
rect -211 19 -207 23
rect -203 20 -202 23
rect -203 19 -100 20
rect -216 16 -100 19
rect -204 12 -200 16
rect -188 12 -184 16
rect -158 12 -154 16
rect -142 12 -138 16
rect -104 12 -100 16
rect -212 -19 -208 8
rect -196 4 -192 8
rect -180 4 -176 8
rect -196 0 -176 4
rect -172 -3 -168 8
rect -150 4 -146 8
rect -134 4 -130 8
rect -150 0 -130 4
rect -124 -3 -120 8
rect -201 -7 -131 -3
rect -124 -7 -100 -3
rect -196 -15 -176 -11
rect -196 -19 -192 -15
rect -180 -19 -176 -15
rect -172 -19 -168 -7
rect -150 -15 -130 -11
rect -150 -19 -146 -15
rect -134 -19 -130 -15
rect -124 -19 -120 -7
rect -93 -19 -89 8
rect -62 -1 -56 37
rect 37 38 190 42
rect -4 27 10 28
rect 33 27 50 31
rect 54 27 66 31
rect 70 27 92 31
rect -4 23 -3 27
rect 1 23 5 27
rect 9 24 10 27
rect 9 23 112 24
rect -4 20 112 23
rect 8 16 12 20
rect 24 16 28 20
rect 54 16 58 20
rect 70 16 74 20
rect 108 16 112 20
rect 0 -1 4 12
rect 16 8 20 12
rect 32 8 36 12
rect 16 4 36 8
rect 40 1 44 12
rect 62 8 66 12
rect 78 8 82 12
rect 62 4 82 8
rect 88 1 92 12
rect -62 -6 4 -1
rect 11 -3 81 1
rect 88 -3 112 1
rect 0 -15 4 -6
rect 16 -11 36 -7
rect 16 -15 20 -11
rect 32 -15 36 -11
rect 40 -15 44 -3
rect 62 -11 82 -7
rect 62 -15 66 -11
rect 78 -15 82 -11
rect 88 -15 92 -3
rect 119 -15 123 12
rect 185 -3 190 38
rect 344 36 348 47
rect 303 25 317 26
rect 340 25 357 29
rect 361 25 373 29
rect 377 25 399 29
rect 303 21 304 25
rect 308 21 312 25
rect 316 22 317 25
rect 316 21 419 22
rect 303 18 419 21
rect 315 14 319 18
rect 331 14 335 18
rect 361 14 365 18
rect 377 14 381 18
rect 415 14 419 18
rect 307 -3 311 10
rect 323 6 327 10
rect 339 6 343 10
rect 323 2 343 6
rect 347 -1 351 10
rect 369 6 373 10
rect 385 6 389 10
rect 369 2 389 6
rect 395 -1 399 10
rect 185 -9 311 -3
rect 318 -5 388 -1
rect 395 -5 419 -1
rect 307 -17 311 -9
rect 323 -13 343 -9
rect 323 -17 327 -13
rect 339 -17 343 -13
rect -204 -35 -200 -23
rect -188 -35 -184 -23
rect -158 -35 -154 -23
rect -142 -35 -138 -23
rect -104 -35 -100 -23
rect 8 -31 12 -19
rect 24 -31 28 -19
rect 54 -31 58 -19
rect 70 -31 74 -19
rect 108 -31 112 -19
rect 347 -17 351 -5
rect 369 -13 389 -9
rect 369 -17 373 -13
rect 385 -17 389 -13
rect 395 -17 399 -5
rect 426 -17 430 10
rect 457 3 462 47
rect 515 29 529 30
rect 552 29 569 33
rect 573 29 585 33
rect 589 29 611 33
rect 515 25 516 29
rect 520 25 524 29
rect 528 26 529 29
rect 528 25 631 26
rect 515 22 631 25
rect 527 18 531 22
rect 543 18 547 22
rect 573 18 577 22
rect 589 18 593 22
rect 627 18 631 22
rect 519 3 523 14
rect 535 10 539 14
rect 551 10 555 14
rect 535 6 555 10
rect 559 3 563 14
rect 581 10 585 14
rect 597 10 601 14
rect 581 6 601 10
rect 607 3 611 14
rect 457 -2 523 3
rect 530 -1 600 3
rect 607 -1 631 3
rect 519 -13 523 -2
rect 535 -9 555 -5
rect 535 -13 539 -9
rect 551 -13 555 -9
rect 559 -13 563 -1
rect 581 -9 601 -5
rect 581 -13 585 -9
rect 597 -13 601 -9
rect 607 -13 611 -1
rect 638 -13 642 14
rect -216 -38 -100 -35
rect -216 -42 -215 -38
rect -211 -42 -207 -38
rect -203 -39 -100 -38
rect -4 -34 112 -31
rect 315 -33 319 -21
rect 331 -33 335 -21
rect 361 -33 365 -21
rect 377 -33 381 -21
rect 415 -33 419 -21
rect 527 -29 531 -17
rect 543 -29 547 -17
rect 573 -29 577 -17
rect 589 -29 593 -17
rect 627 -29 631 -17
rect -4 -38 -3 -34
rect 1 -38 5 -34
rect 9 -35 112 -34
rect 9 -38 10 -35
rect -4 -39 10 -38
rect 303 -36 419 -33
rect -203 -42 -202 -39
rect 303 -40 304 -36
rect 308 -40 312 -36
rect 316 -37 419 -36
rect 515 -32 631 -29
rect 515 -36 516 -32
rect 520 -36 524 -32
rect 528 -33 631 -32
rect 528 -36 529 -33
rect 515 -37 529 -36
rect 316 -40 317 -37
rect 303 -41 317 -40
rect -216 -43 -202 -42
<< labels >>
rlabel metal1 -1 22 -1 22 1 VDD
rlabel metal1 11 -33 11 -33 1 Gnd
rlabel metal1 -213 18 -213 18 1 VDD
rlabel metal1 -201 -37 -201 -37 1 Gnd
rlabel metal1 518 24 518 24 1 VDD
rlabel metal1 640 -1 640 -1 1 Sum0
rlabel metal1 530 -31 530 -31 1 Gnd
rlabel metal1 306 20 306 20 1 VDD
rlabel metal1 318 -35 318 -35 1 Gnd
rlabel metal1 428 -5 428 -5 1 Sum1
rlabel polycontact 558 38 558 38 1 cin0
rlabel metal1 520 1 520 1 1 cout0
rlabel polycontact 337 27 337 27 1 b1
rlabel polycontact 329 27 329 27 1 a1
rlabel metal1 308 -3 308 -3 1 cout1
rlabel polycontact 541 31 541 31 1 a1
rlabel polycontact 549 31 549 31 1 b1
rlabel metal1 121 -3 121 -3 1 sum2
rlabel polycontact 30 29 30 29 1 b2
rlabel polycontact 22 29 22 29 1 a1
rlabel metal1 1 -1 1 -1 1 cout2
rlabel metal1 -91 -8 -91 -8 1 sum3
rlabel polycontact -182 25 -182 25 1 b3
rlabel polycontact -190 25 -190 25 1 a3
rlabel metal1 -211 -5 -211 -5 1 cout3
<< end >>
