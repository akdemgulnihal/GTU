magic
tech scmos
timestamp 1699549236
<< nwell >>
rect -3 -7 22 21
<< ntransistor >>
rect 9 -20 11 -16
<< ptransistor >>
rect 9 0 11 8
<< ndiffusion >>
rect 8 -20 9 -16
rect 11 -20 12 -16
<< pdiffusion >>
rect 8 4 9 8
rect 4 0 9 4
rect 11 4 16 8
rect 11 0 12 4
<< ndcontact >>
rect 4 -20 8 -16
rect 12 -20 16 -16
<< pdcontact >>
rect 4 4 8 8
rect 12 0 16 4
<< psubstratepcontact >>
rect 1 -29 5 -25
rect 15 -29 19 -25
<< nsubstratencontact >>
rect 1 13 5 17
rect 15 13 19 17
<< polysilicon >>
rect 9 8 11 11
rect 9 -6 11 0
rect 7 -10 11 -6
rect 9 -16 11 -10
rect 9 -23 11 -20
<< polycontact >>
rect 3 -10 7 -6
<< metal1 >>
rect 0 17 20 18
rect 0 13 1 17
rect 5 13 15 17
rect 19 13 20 17
rect 0 12 20 13
rect 4 8 8 12
rect -1 -10 3 -6
rect 12 -16 16 0
rect 4 -24 8 -20
rect 0 -25 20 -24
rect 0 -29 1 -25
rect 5 -29 15 -25
rect 19 -29 20 -25
rect 0 -30 20 -29
<< labels >>
rlabel metal1 6 -27 6 -27 1 gnd
rlabel metal1 -1 -8 -1 -8 3 input
rlabel metal1 16 -8 16 -8 7 output
rlabel metal1 6 15 6 15 5 vdd
<< end >>
